module FOUR_4bit( output [3:0] out );
  assign out = 4'b0100;
endmodule
