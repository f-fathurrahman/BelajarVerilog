module main;
  initial
  begin
    $display("Hello from ffr");
    $finish;
  end
endmodule

