module test1( in1, out1 );
  input in1;
  output out1;
  
  assign out1 = in1;
endmodule;
