module THREE_4bit( output [3:0] out );
  assign out = 4'b0011;
endmodule 
