module tes_led8( output [7:0] led);

  assign led = 8'b0100_0000;

endmodule
