module HIGH(output out);
  assign out = 1;
endmodule
