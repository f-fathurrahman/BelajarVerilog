module LOW( output out);
  assign out = 0;
endmodule
