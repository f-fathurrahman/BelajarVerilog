module TWO_4bit( output [3:0] out );
  assign out = 4'b0010;
endmodule
